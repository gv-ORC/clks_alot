module top (
    // input  common_p::clk_dom_s sys_dom_i, //! Use the init/config handshake



    output clks_alot_p::clock_status_s recover_status_o, // Recovery

    output clks_alot_p::generated_events_s actual_clks_o,    // Recovery
    output clks_alot_p::generated_events_s expected_clks_o,  // Generation
    output clks_alot_p::generated_events_s preemetive_clks_o // Generation
);

// Recovery

// 

endmodule : top
