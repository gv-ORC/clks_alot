/*
1. Recover Events
2. Send Events to the appropriate one (of two) `rate_recovery` modules
3. Forward Events and Rates to generation system
*/
